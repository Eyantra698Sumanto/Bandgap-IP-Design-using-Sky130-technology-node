* SPICE3 file created from starternfet.ext - technology: sky130A

.subckt starternfet net6 gnd
X0 a_88_252# a_88_252# gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=7e+06u
X1 net6 net6 a_88_252# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=7e+06u
C0 net6 gnd 2.30fF
C1 a_88_252# gnd 2.69fF
.ends
